`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// zero_extend_12_to_16.sv
//////////////////////////////////////////////////////////////////////////////////

module zero_extend_12_to_16(
    input  logic [11:0] in12,
    output logic [15:0] out16
);
    assign out16 = {4'd0, in12};
endmodule
