module averager_pwm
    #(parameter int
        power = 8, // 2**power samples, default is 2**8 = 256 samples
        N     = 12 // # of bits to take the average of
    )
    (
        input  logic          clk,
        input  logic          reset,
        input  logic          EN,
        input  logic [N-1:0]  Din,   // input to averager
        output logic [N-1:0]  Q      // N-bit moving average
    );

    // Storage for last 2**power samples (1-based indexing to match your other code)
    logic [N-1:0] REG_ARRAY [2**power:1];

    // Running sum of window (needs N + power bits)
    logic [power+N-1:0] sum;

    // Average = sum / 2**power  -> just take upper bits
    assign Q = sum[power+N-1:power];

    always_ff @(posedge clk) begin
        if (reset) begin
            sum <= '0;
            for (int j = 1; j <= 2**power; j++) begin
                REG_ARRAY[j] <= '0;
            end
        end
        else if (EN) begin
            // Sliding-window: remove oldest, add newest
            sum <= sum + Din - REG_ARRAY[2**power];

            // Shift register contents "down"
            for (int j = 2**power; j > 1; j--) begin
                REG_ARRAY[j] <= REG_ARRAY[j-1];
            end

            // Insert newest sample at the front
            REG_ARRAY[1] <= Din;
        end
    end

endmodule
