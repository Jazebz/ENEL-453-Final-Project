`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// zero_extend_8_to_16.sv
//////////////////////////////////////////////////////////////////////////////////

module zero_extend_8_to_16(
    input  logic [7:0]  in8,
    output logic [15:0] out16
);
    assign out16 = {8'd0, in8};
endmodule
